// to learn more about VGA control design, type:
// https://www.intel.com/content/dam/support/us/en/programmable/support-resources/fpga-wiki/asset03/basic-vga-controller-design-example.pdf

module vga(
		input vgaclk,           //input pixel clock: how fast should this be? // megaclock / 2
		input rst,              //synchronous reset
		output hsync,			//horizontal sync out
		output vsync,			//vertical sync out
		output reg [3:0] red,	//red vga output
		output reg [3:0] green, //green vga output
		output reg [3:0] blue	//blue vga output
   );
// VGA: 480 X 640 module
// VGA protocol: 
	
	// refresh rate = 60Hz
	// TODO: Video protocol constants
   // You can find these described in the VGA specification for 640x480
	localparam HPIXELS = 639;  // horizontal pixels per line
	localparam HBP = HPIXELS + 16; 	// end of horizontal back porch
	localparam HFP = HBP + 96; 	    // hsync pulse length
	localparam TOTALH = HFP + 48; 	    // beginning of horizontal front porch
	
	localparam VLINES = 479;   // scanlines per frame (aka the # of vertical pixels)
	localparam VBP = VLINES + 10; 		// end of vertical back porch
	localparam VFP = VBP + 2; 	    // beginning of vertical front porch
	localparam TOTALV = VFP + 33; 	// vsync pulse length
	
	localparam rr = 60; // refresh rate
	// registers for storing the horizontal & vertical counters
	reg [9:0] hc = 0;
	reg [9:0] vc = 0;
	reg de = 0; // LOW if blanking interval, HIGH if printing
	reg [18:0] counter = 19'h0;
	// doesn't work unless in testbench // reg[3:0] seed = 4'hF; // random number generator seed
	// doesn't work unless in testbench // reg[31:0] randval; // random value generated by $urandom()
	
    //Counter block: change hc and vc correspondingly to the current state.
	always @(posedge vgaclk) begin
		 //reset condition
		if (rst == 1)
		begin
			hc<=0;
			vc<=0;
			counter<=0;
		end
		else if (hc >= 799)
		begin
			hc<=0;
			vc<=vc+1;
			if (vc >= 524) begin
				hc<=0;
				vc<=0;
				counter<=0;
			end 
		end
		else begin
			//TODO: Implement logic to move counters properly!
			hc<=hc+1;
			counter<=counter+1;
		end
	end

	assign hsync = ~((hc > HBP) && (hc <= HFP)); 
	assign vsync = ~((vc > VBP) && (vc <= VFP));
	
	//RGB output block: set red, green, blue outputs here.
	always@(posedge vgaclk)
	begin
		// check if we're within vertical active video range
		if ( ( 300<hc && hc<340) && ( 200<vc && vc<280 ) )  // the screen is 640 * 480 ==> divide by 8 (80 * 400)
		begin
			//TODO: draw something!
			red <= 4'hF;
			green <= 4'hF;
			blue <= 4'h0;
		end
		else if( (0 <= hc && hc < 80) && (0 <= vc && vc < 400))
		begin
			red <= 4'hF;
			green <= 4'h0;
			blue <= 4'h0;
		end
		else if( (80<=hc && hc<160) && (0<=vc && vc<400))
		begin
			red <= 4'hF;
			green <= 4'h8;
			blue <= 4'h0;
		end
		else if( (160<= hc && hc < 240) && (0<=vc && vc<400))
		begin
			red <= 4'hF;
			green <= 4'hF;
			blue <= 4'h0;
		end
		else if( (240<=hc && hc<320) && (0<=vc && vc<400))
		begin
			red <= 4'h0;
			green <= 4'hF;
			blue <= 4'h0;
		end
		else if( (320<= hc && hc < 400) && (0<=vc && vc<400))
		begin
			red <= 4'h0;
			green <= 4'hF;
			blue <= 4'h8;
		end
		else if( (400<=hc && hc<480) && (0<=vc && vc<400))
		begin
			red <= 4'h0;
			green <= 4'hF;
			blue <= 4'hF;
		end
		else if( (480<= hc && hc < 560) && (0<=vc && vc<400))
		begin
			red <= 4'h0;
			green <= 4'h8;
			blue <= 4'hF;
		end
		else if( (560<=hc && hc<640) && (0<=vc && vc<400))
		begin
			red <= 4'h0;
			green <= 4'h0;
			blue <= 4'hF;
		end
		else begin
			//TODO: we're not in active video range, what do we do?
			// black screen
			red <= 4'h0;
			green <= 4'h0;
			blue <= 4'h0;
		end
	end

endmodule
