module butteryfly_16();

endmodule